'default_nettype none
